module testbench;
  reg a_tb; reg b_tb; wire y_tb;
  XOR_1 uut(a_tb,b_tb,y_tb);
  initial begin 
    $dumpfile("dump.vcd");
    $dumpvars(0, testbench);
  end
  
  initial
    begin
      $monitor($time,"a_tb=%b, b_tb=%b, y_tb=%b",a_tb,b_tb,y_tb);
      
      #5 a_tb=0; b_tb=0;
      #5 a_tb=0; b_tb=1;
      #5 a_tb=1; b_tb=0;
      #5 a_tb=1; b_tb=1;
      #5 $finish;
    end
endmodule
